`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   00:06:44 06/05/2021
// Design Name:   parking_meter
// Module Name:   /home/ise/xilinx/Proj4/Proj4/testbench_305330193.v
// Project Name:  Proj4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: parking_meter
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testbench_305330193;

	reg add1;
	reg add2;
	reg add3;
	reg add4;
	reg rst1;
	reg rst2;
	reg clk;
	reg rst;
	// Outputs
	wire [6:0] led_seg;
	wire a1;
   wire a2;
   wire a3;
   wire a4;
	wire [3:0] val1;
	wire [3:0] val2;
	wire [3:0] val3;
	wire [3:0] val4;

	// Instantiate the Unit Under Test (UUT)
	parking_meter uut (
		.add1(add1), 
		.add2(add2), 
		.add3(add3), 
		.add4(add4), 
		.rst1(rst1), 
		.rst2(rst2), 
		.clk(clk), 
		.rst(rst), 
		.led_seg(led_seg),
		.a1(a1),
		.a2(a2),
		.a3(a3),
		.a4(a4),
		.val1(val1),
		.val2(val2),
		.val3(val3),
		.val4(val4)
	);

	initial begin
		// Initialize Inputs
		add1 = 0;
		add2 = 0;
		add3 = 0;
		add4 = 0;
		rst1 = 0;
		rst2 = 0;
		clk = 0;
		rst = 0;
		
     //see if add inputs work fine
		rst = 1;
		#5000000
		rst = 0;
		#10000000
		add1 = 1;
		#1000000000
		add1 = 0;
		#1000000000
		add2 = 1;
		#1000000000
		add2 = 0;
		#1000000000
		add3 = 1;
		#1000000000
		add3 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		//wait 10s
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		rst1 = 1;
		#100000000
		rst1 = 0;
		//wait 10s
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		//reset it to 150 seconds
		rst2 = 1;
		#50
		rst2 = 0;
		//wait 5 sec
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		//there will be bunch of add4 to hit the 9999 mark and check if it stays 9999 when add4 at 9999 sec
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000 
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		#1000000000
		add4 = 1;
		#1000000000
		add4 = 0;
		//wait 10 s to see the decrement and flashing when > 180
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		//see the reset works
		rst = 1;
		#1000000000
		rst = 0;
		//check the flashing at 0 sec (1s with 50% duty cycle)
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		//change the time to 150
		rst2 = 1;
		#1000000000
		rst2 = 0;
		//and increment it by 60
		#1000000000
		add1 = 1;
		#1000000000
		add1 = 0;
		//seconds > 180 so always flash
		//40 seconds of wait --> flashing should transition to 2s 50% duty cycle
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		//reset to 16 and watch it count down
		rst1 = 1;
		#1000000000
		rst1 =0;
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		#1000000000
		$stop;
	end
	always clk = #5000000 ~clk;
      
endmodule

